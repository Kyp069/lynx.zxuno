//-------------------------------------------------------------------------------------------------
module audio
//-------------------------------------------------------------------------------------------------
(
	input  wire      clock,
	input  wire      reset,
	input  wire      ear,
	input  wire[5:0] dac,
	output wire[1:0] audio
);
//-------------------------------------------------------------------------------------------------

reg source;
always @(posedge clock) source <= ~source;

wire[5:0] mix = source ? {6{ear}} : dac;

//-------------------------------------------------------------------------------------------------

dac #(.MSBI(5)) Dac
(
	.clock(clock  ),
	.reset(reset  ),
	.di   (mix    ),
	.do   (dacDo  )
);

assign audio = {2{dacDo}};

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
