//-------------------------------------------------------------------------------------------------
module spr
//-------------------------------------------------------------------------------------------------
#
(
	parameter DW = 8,
	parameter AW = 14
)
(
	input  wire         clock,
	input  wire         ce,
	input  wire         we,
	input  wire[   7:0] di,
	output reg [   7:0] do,
	input  wire[AW-1:0] a
);
//-------------------------------------------------------------------------------------------------

reg[7:0] d[(2**AW)-1:0];

always @(posedge clock) if(ce) if(!we) d[a] <= di; else do <= d[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
